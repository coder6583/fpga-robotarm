`default_nettype none

module Jacobian
    ();
endmodule : Jacobian
